// Synchronous FIFO

module sync (
    
);

endmodule //sync